module vgama

import gg

const keys = {
	// Direction keys -> 'd' class (direction)
	gg.KeyCode.invalid:       '  '
	gg.KeyCode.up:            'au'
	gg.KeyCode.down:          'ad'
	gg.KeyCode.left:          'al'
	gg.KeyCode.right:         'ar'
	// Special keys -> 's' class (special/control)
	gg.KeyCode.escape:        'sx'
	gg.KeyCode.insert:        'si'
	gg.KeyCode.delete:        'sd'
	gg.KeyCode.home:          'sh'
	gg.KeyCode.end:           'sn'
	gg.KeyCode.page_up:       'su'
	gg.KeyCode.page_down:     'sp'
	// Modifiers -> 'm' class (modifiers)
	gg.KeyCode.left_shift:    'ms'
	gg.KeyCode.right_shift:   'ms'
	gg.KeyCode.left_control:  'mc'
	gg.KeyCode.right_control: 'mc'
	gg.KeyCode.left_alt:      'ma'
	gg.KeyCode.right_alt:     'ma'
	gg.KeyCode.left_super:    'mS'
	gg.KeyCode.right_super:   'mS'
	gg.KeyCode.caps_lock:     'mC'
	// Character keys -> 'c' class (character)
	gg.KeyCode.a:             'ca'
	gg.KeyCode.b:             'cb'
	gg.KeyCode.c:             'cc'
	gg.KeyCode.d:             'cd'
	gg.KeyCode.e:             'ce'
	gg.KeyCode.f:             'cf'
	gg.KeyCode.g:             'cg'
	gg.KeyCode.h:             'ch'
	gg.KeyCode.i:             'ci'
	gg.KeyCode.j:             'cj'
	gg.KeyCode.k:             'ck'
	gg.KeyCode.l:             'cl'
	gg.KeyCode.m:             'cm'
	gg.KeyCode.n:             'cn'
	gg.KeyCode.o:             'co'
	gg.KeyCode.p:             'cp'
	gg.KeyCode.q:             'cq'
	gg.KeyCode.r:             'cr'
	gg.KeyCode.s:             'cs'
	gg.KeyCode.t:             'ct'
	gg.KeyCode.u:             'cu'
	gg.KeyCode.v:             'cv'
	gg.KeyCode.w:             'cw'
	gg.KeyCode.x:             'cx'
	gg.KeyCode.y:             'cy'
	gg.KeyCode.z:             'cz'
	// Digits
	gg.KeyCode._0:            'c0'
	gg.KeyCode._1:            'c1'
	gg.KeyCode._2:            'c2'
	gg.KeyCode._3:            'c3'
	gg.KeyCode._4:            'c4'
	gg.KeyCode._5:            'c5'
	gg.KeyCode._6:            'c6'
	gg.KeyCode._7:            'c7'
	gg.KeyCode._8:            'c8'
	gg.KeyCode._9:            'c9'
	// Whitespace and punctuation
	gg.KeyCode.space:         'c '
	gg.KeyCode.tab:           'c\t'
	gg.KeyCode.enter:         'c\n'
	gg.KeyCode.comma:         'c,'
	gg.KeyCode.period:        'c.'
	gg.KeyCode.slash:         'c/'
	gg.KeyCode.semicolon:     'c;'
	gg.KeyCode.apostrophe:    "c'"
	gg.KeyCode.backslash:     'c\\'
	gg.KeyCode.left_bracket:  'c['
	gg.KeyCode.right_bracket: 'c]'
	gg.KeyCode.minus:         'c-'
	gg.KeyCode.equal:         'c='
	// Function keys -> 'f' class (function)
	gg.KeyCode.f1:            'f1'
	gg.KeyCode.f2:            'f2'
	gg.KeyCode.f3:            'f3'
	gg.KeyCode.f4:            'f4'
	gg.KeyCode.f5:            'f5'
	gg.KeyCode.f6:            'f6'
	gg.KeyCode.f7:            'f7'
	gg.KeyCode.f8:            'f8'
	gg.KeyCode.f9:            'f9'
	gg.KeyCode.f10:           'fa'
	gg.KeyCode.f11:           'fb'
	gg.KeyCode.f12:           'fc'
}
