module main

import gg

fn c_redimension(x f64, y f64, w f64, h f64) (f32, f32, f32, f32) {
	return f32((x + 1) * width), f32((y + 1) * height), f32(w * height), f32(h * height)
}

fn c_color(r u8, g u8, b u8, _ u8) gg.Color {
	return gg.rgb(r, g, b)
}
