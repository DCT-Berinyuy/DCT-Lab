module vgama

interface Compiler {
}
